*
* MODELO SPICE
*

* para guardar as correntes
.options savecurrents


* alimentacao
Vcc vcc 0 5.0
Vee vee 0 -5.0
I1 ve 0 200u

* fonte de entrada
Vin 1 0 0.0 ac 1.0 sin(0 .1 100k)

Rs 1 vb1 10k
Rc1 vcc vc1 38k
Rc2 vcc vc2 38k
Rl vc3 0 2k
Cc vx vb2 1

R1 vb2 0 1k
R2 vx ve3 10k
Re vcc ve3 1k


Q1 vc1 vb1 ve Nmodel
Q2 vc2 vb2 ve Nmodel
Q3 vc3 vb3 ve3 Pmodel


.model Nmodel NPN(Bf=400, CJE=12pF, CJC=2pF)
.model Pmodel NPN(Bf=600, CJE=12pF, CJC=2pF)

.end


*PFR
*op
*print @q1[ic]

* analise no tempo
*tran 1e-5 10e-3

*análise na frequência
*ac dec 10 10 100MEG
*plot db(v(coll))
*plot vp(coll)

*impedancia de entrada
*print v(2)[40]/abs(v(2)[40]-v(1)[40])*1000