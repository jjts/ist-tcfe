*
* MODELO SPICE
* Retificador de meia onda com deslocamento de nivel DC
*


* subcircuito do ampop
.subckt opamp plus minus out
*
r1 plus minus 300k
a1 %vd (plus minus) outint lim
.model lim limit (out_lower_limit = -12 out_upper_limit = 12
+ fraction = true limit_range = 0.2 gain=300e3)
r3 outint out 50.0
r2 out 0 1e12
*
.ends opamp
*


* para guardar as correntes
.options savecurrents

*
*
*
* fonte de entrada
Vin i 0 sin(6 2 1000)
*
*
*
*

* passa-alto ordem 1 a entrada 
Ci i 1 100u
Rhp 1 0 10k


* ampop
xampop 1 2 2 opamp

* detector de envolvente (rectificador + passa-baixo)
D0 2 o DMOD
Co o 0 100u
Ro o 0 10k


* modelo do diodo

.model DMOD D (bv=50 is=1e-13 n=1.05)
.model Da1N4004 D (IS=18.8n RS=0 BV=400 IBV=5.00u M=0.333 N=2)

.end


* COMMANDS


* analise no tempo
* tran 1e-5 1
*plot v(i) v(o)


