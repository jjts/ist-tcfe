*
* MODELO SPICE
* Amp BJT Realimentado
*

* para guardar as correntes
.options savecurrents


* alimentacao
Vcc vcc 0 10.0

* fonte de entrada
Vin 1 0 0.0 ac 1.0 sin(0 .1 100k)

Rs 1 2 1k

* condensador de acoplamento à entrada
Cb 2 base 1uF

Rf coll base 50k

Q1 coll base emit P2model

Rc vcc coll 300

Re emit 0 100

Ce emit 0 10uF

.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)

.end


*PFR
*op
*print @q1[ic]

* analise no tempo
*tran 1e-5 10e-3

*análise na frequência
*ac dec 10 10 100MEG
*plot db(v(coll))
*plot vp(coll)

*impedancia de entrada
*print v(2)[40]/abs(v(2)[40]-v(1)[40])*1000