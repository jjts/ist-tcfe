*
* MODELO SPICE
* Filtro de Rauch
*


* subcircuito do ampop
.subckt opamp plus minus out
*
r1 plus minus 300k
a1 %vd (plus minus) outint lim
.model lim limit (out_lower_limit = -12 out_upper_limit = 12
+ fraction = true limit_range = 0.2 gain=300e3)
r3 outint out 50.0
r2 out 0 1e12
*
.ends opamp
*


* para guardar as correntes
.options savecurrents

*
*
*
* fonte de entrada
Vin i 0 ac 1.0 sin(0 1 1000)
*
*
*
*

* ampop
xampop 0 vminus o opamp

R1 i 1 11.251k
C2 1 0  3n
R3 1 vminus  11.251k
R4 1 o  11.251k
C5 vminus o 667p

.end


* comandos

*análise na frequência
*ac dec 10 10 100MEG
*plot vdb(o)
*plot phase(o)


